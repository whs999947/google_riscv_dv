module top;
initial begin
  $display("hello sv");
end
endmodule
